library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--Asteroid Sprite Table
entity asteroid_sprite_table is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(63 downto 0)
   );
end asteroid_sprite_table;

architecture arch of asteroid_sprite_table is
   
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=64;
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
   
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
        
   -- ROM definition
   constant ROM: rom_type:=( 
     -- code x00
   "0000000000000000000000000000000000001111110000000000000000000000", -- 00
   "0000000000000000000000000000000000010000001000000000000000000000", -- 01
   "0000000000000000000000000000000000100000000100000000000000000000", -- 02
   "0000000000000000000000000000000001000000000010000000000000000000", -- 03
   "0000000000000000000000000000000010000000000001000000000000000000", -- 04
   "0000000000000000000000000000000100000000000000100000000000000000", -- 05
   "0000000000000000000000000000001000000000000000010000000000000000", -- 06
   "0000000000000000000000000011111000000000000000001000000000000000", -- 07
   "0000000000000000000000000100000000000000000000000100000000000000", -- 08
   "0000000000000000000000001000000000000000000000000011111111000000", -- 09
   "0000000000000000000000010000000000000000000000000000000000100000", -- 0a
   "0000000000000000000000100000000000000000000000000000000000010000", -- 0b
   "0000000000000000000001000000000000000000000000000000000000001000", -- 0c
   "0000000000000000000010000000000000000000000000000000000000000100", -- 0d
   "0000000000000000000100000000000000000000000000000000000000000010", -- 0e
   "0000000000000000001000000000000000000000000000000000000000000010", -- 0f
   "0000000000000000010000000000000000000000000000000000000000000010", -- 10
   "0000000000000000100000000000000000000000000000000000000000000010", -- 11
   "0000000000000000100000000000000000000000000000000000000000000010", -- 12
   "0000000000000000100000000000000000000000000000000000000000000010", -- 13
   "0000000000000000100000000000000000000000000000000000000000000100", -- 14
   "0000000000000000100000000000000000000000000000000000000000001000", -- 15
   "0000000000000000100000000000000000000000000000000000000000010000", -- 16
   "0000000000000000100000000000000000000000000000000000000000100000", -- 17
   "0000000000000000100000000000000000000000000000000000000001000000", -- 18
   "0000000000000000100000000000000000000000000000000000000010000000", -- 19
   "0000000000000000010000000000000000000000000000000000000100000000", -- 1a
   "0000000000000000001000000000000000000000000000000000001000000000", -- 1b
   "0000000000000000000100000000000000000000000000000000010000000000", -- 1c
   "0000000000000000000010000000000000000000000000000000010000000000", -- 1d
   "0000000000000000000001000000000000000000000000000000010000000000", -- 1e
   "0000000000000000000000100000000000000000000000000000001000000000", -- 1f
   "0000000000000000000000010000000000000000000000000000000100000000", -- 20
   "0000000000000000000000100000000000000000000000000000000010000000", -- 21
   "0000000000000000000001000000000000000000000000000000000001000000", -- 22
   "0000000000000000000010000000000000000000000000000000000000100000", -- 23
   "0000000000000000000100000000000000000000000000000000000000010000", -- 24
   "0000000000000000001000000000000000000000000000000000000000001000", -- 25
   "0000000000000000010000000000000000000000000000000000000000001000", -- 26
   "0000000000000000100000000000000000000000000000000000000000001000", -- 27
   "0000000000000000100000000000000000000000000000000000000000001000", -- 28
   "0000000000000000100000000000000000000000000000000000000000001000", -- 29
   "0000000000000000010000000000000000000000000000000000000000001000", -- 2a
   "0000000000000000001000000000000000000000000000000000000000001000", -- 2b
   "0000000000000000000100000000000000000000000000000000000000001000", -- 2c
   "0000000000000000000010000000000000000000000000000000000000001000", -- 2d
   "0000000000000000000001000000000000000000000000000000000000001000", -- 2e
   "0000000000000000000000100000000000000000000000000000000000010000", -- 2f
   "0000000000000000000000010000000000000000000000000000000000100000", -- 30
   "0000000000000000000000010000000000000000000000000000000001000000", -- 31
   "0000000000000000000000010000000000000000000000000000000010000000", -- 32
   "0000000000000000000000010000000000000000000000000000000100000000", -- 33
   "0000000000000000000000010000000000000000000000000000001000000000", -- 34
   "0000000000000000000000010000000000000000000000000000010000000000", -- 35
   "0000000000000000000000010000000000000000000000000000100000000000", -- 36
   "0000000000000000000000010000000000000000000000000001000000000000", -- 37
   "0000000000000000000000010000000000000001111111111110000000000000", -- 38
   "0000000000000000000000010000000000000010000000000000000000000000", -- 39
   "0000000000000000000000001000000000000100000000000000000000000000", -- 3a
   "0000000000000000000000000100000000001000000000000000000000000000", -- 3b
   "0000000000000000000000000011111111110000000000000000000000000000", -- 3c
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3d
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3e
   "0000000000000000000000000000000000000000000000000000000000000000",  -- 3f
     -- code x01
   "0000000000000000000000000000000000000000000000000000000000000000", -- 00
   "0000000000000000000000001111111111111100000000000000000000000000", -- 01
   "0000000000000000000000010000000000000010000000000000000000000000", -- 02
   "0000000000000000000000100000000000000001000000000000000000000000", -- 03
   "0000000000000000000001000000000000000000100000000000000000000000", -- 04
   "0000000000000000000010000000000000000000011111111100000000000000", -- 05
   "0000000000000000000100000000000000000000000000000011000000000000", -- 06
   "0000000000011111111000000000000000000000000000000000110000000000", -- 07
   "0000000000100000000000000000000000000000000000000000001100000000", -- 08
   "0000000001000000000000000000000000000000000000000000000011000000", -- 09
   "0000000010000000000000000000000000000000000000000000000000110000", -- 0a
   "0000000100000000000000000000000000000000000000000000000000001000", -- 0b
   "0000001000000000000000000000000000000000000000000000000000000100", -- 0c
   "0000010000000000000000000000000000000000000000000000000000000100", -- 0d
   "0000010000000000000000000000000000000000000000000000000000000100", -- 0e
   "0000010000000000000000000000000000000000000000000000000000000100", -- 0f
   "0000001000000000000000000000000000000000000000000000000000000100", -- 10
   "0000000100000000000000000000000000000000000000000000000000000100", -- 11
   "0000000010000000000000000000000000000000000000000000000000001000", -- 12
   "0000000010000000000000000000000000000000000000000000000000010000", -- 13
   "0000000010000000000000000000000000000000000000000000000000100000", -- 14
   "0000000001100000000000000000000000000000000000000000000001000000", -- 15
   "0000000000011000000000000000000000000000000000000000000010000000", -- 16
   "0000000000000110000000000000000000000000000000000000000100000000", -- 17
   "0000000000000001100000000000000000000000000000000000001000000000", -- 18
   "0000000000000000100000000000000000000000000000000000001000000000", -- 19
   "0000000000000000100000000000000000000000000000000000001000000000", -- 1a
   "0000000000000001000000000000000000000000000000000000001000000000", -- 1b
   "0000000000000010000000000000000000000000000000000000001000000000", -- 1c
   "0000000000000100000000000000000000000000000000000000001000000000", -- 1d
   "0000000000001000000000000000000000000000000000000000001000000000", -- 1e
   "0000000000010000000000000000000000000000000000000000010000000000", -- 1f
   "0000000000100000000000000000000000000000000000000000100000000000", -- 20
   "0000000001000000000000000000000000000000000000000001000000000000", -- 21
   "0000000001000000000000000000000000000000000000000010000000000000", -- 22
   "0000000001000000000000000000000000000000000000000100000000000000", -- 23
   "0000000000100000000000000000000001000000000000001000000000000000", -- 24
   "0000000000010000000000000000000010100000000000010000000000000000", -- 25
   "0000000000001000000000000000000100010000000000100000000000000000", -- 26
   "0000000000000100000000000000001000001000000001000000000000000000", -- 27
   "0000000000000010000000000000010000000111111110000000000000000000", -- 28
   "0000000000000001000000000000100000000000000000000000000000000000", -- 29
   "0000000000000000100000000001000000000000000000000000000000000000", -- 2a
   "0000000000000000011111111110000000000000000000000000000000000000", -- 2b
   "0000000000000000000000000000000000000000000000000000000000000000", -- 2c
   "0000000000000000000000000000000000000000000000000000000000000000", -- 2d
   "0000000000000000000000000000000000000000000000000000000000000000", -- 2e
   "0000000000000000000000000000000000000000000000000000000000000000", -- 2f
   "0000000000000000000000000000000000000000000000000000000000000000", -- 30
   "0000000000000000000000000000000000000000000000000000000000000000", -- 31
   "0000000000000000000000000000000000000000000000000000000000000000", -- 32
   "0000000000000000000000000000000000000000000000000000000000000000", -- 33
   "0000000000000000000000000000000000000000000000000000000000000000", -- 34
   "0000000000000000000000000000000000000000000000000000000000000000", -- 35
   "0000000000000000000000000000000000000000000000000000000000000000", -- 36
   "0000000000000000000000000000000000000000000000000000000000000000", -- 37
   "0000000000000000000000000000000000000000000000000000000000000000", -- 38
   "0000000000000000000000000000000000000000000000000000000000000000", -- 39
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3a
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3b
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3c
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3d
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3e
   "0000000000000000000000000000000000000000000000000000000000000000",  -- 3f
      -- code x02                                        
   "0000000000000000000000000000000000000000000000000000000000000000", -- 00
   "0000000000000000000000000000000000000000000000000000000000000000", -- 01
   "0000000000000000000000000000000000000000000000000000000000000000", -- 02
   "0000000000000000000000000000000000000000000000000000000000000000", -- 03
   "0000000000000000000000000000000000000000000000000000000000000000", -- 04
   "0000000000000000000000000000000000000000000000000000000000000000", -- 05
   "0000000000000000000000000000000000000000000000000000000000000000", -- 06
   "0000000000000000000000000000000000000000000000000000000000000000", -- 07
   "0000000000000000000000000000000000000000000000000000000000000000", -- 08
   "0000000000000000000000000000000000000000000000000000000000000000", -- 09
   "0000000000000000100000000000000000000000000000001000000000000000", -- 0a
   "0000000000000000100000000000000000000000000000001000000000000000", -- 0b
   "0000000000000111111000000000000000000000000001111110000000000000", -- 0c
   "0000000000001111111100000000000000000000000011111111000000000000", -- 0d
   "0000000000000111111000000000000000000000000001111110000000000000", -- 0e
   "0000000000000000100000000000000000000000000000001000000000000000", -- 0f
   "0000000000000000100000000000000000000000000000001000000000000000", -- 10
   "0000000000000000000000000000000000000000000000000000000000000000", -- 11
   "0000000000000000000000000000000000000000000000000000000000000000", -- 12
   "0000000000000000000000000000000000000000000000000000000000000000", -- 13
   "0000000000000000000000000000000000000000000000000000000000000000", -- 14
   "0000000000000000000000000000000000000000000000000000000000000000", -- 15
   "0000000000000000000000000000000000000000000000000000000000000000", -- 16
   "0000000000000000000000000000000000000000000000000000000000000000", -- 17
   "0000000000000000000000000000000000000000000000000000000000000000", -- 18
   "0000000000000000000000000000000000000000000000000000000000000000", -- 19
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1a
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1b
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1c
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1d
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1e
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1f
   "0000000000000000000000000000000000000000000000000000000000000000", -- 20
   "0000000000000000000000000000000000000000000000000000000000000000", -- 21
   "0000000000000000000000000000000000000000000000000000000000000000", -- 22
   "0000000000000000000000000000000000000000000000000000000000000000", -- 23
   "0000000000000000000000000000000000000000000000000000000000000000", -- 24
   "0000000000000000000000000000000000000000000000000000000000000000", -- 25
   "0000000000000000000000000000000000000000000000000000000000000000", -- 26
   "0000000000000000000000000000000000000000000000000000000000000000", -- 27
   "0000000000000000000000000000000000000000000000000000000000000000", -- 28
   "0000000000000000000000000000000000000000000000000000000000000000", -- 29
   "0000000000000000100000000000000000000000000000001000000000000000", -- 2a
   "0000000000000000100000000000000000000000000000001000000000000000", -- 2b
   "0000000000000111111000000000000000000000000001111110000000000000", -- 2c
   "0000000000001111111100000000000000000000000011111111000000000000", -- 2d
   "0000000000000111111000000000000000000000000001111110000000000000", -- 2e
   "0000000000000000100000000000000000000000000000001000000000000000", -- 2f
   "0000000000000000100000000000000000000000000000001000000000000000", -- 30
   "0000000000000000000000000000000000000000000000000000000000000000", -- 31
   "0000000000000000000000000000000000000000000000000000000000000000", -- 32
   "0000000000000000000000000000000000000000000000000000000000000000", -- 33
   "0000000000000000000000000000000000000000000000000000000000000000", -- 34
   "0000000000000000000000000000000000000000000000000000000000000000", -- 35
   "0000000000000000000000000000000000000000000000000000000000000000", -- 36
   "0000000000000000000000000000000000000000000000000000000000000000", -- 37
   "0000000000000000000000000000000000000000000000000000000000000000", -- 38
   "0000000000000000000000000000000000000000000000000000000000000000", -- 39
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3a
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3b
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3c
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3d
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3e
   "0000000000000000000000000000000000000000000000000000000000000000",  -- 3f
      -- code x03
   "0000000000000000000000000000000000000000000000000000000000000000", -- 00
   "0000000000000000000000000000000000000000000000000000000000000000", -- 01
   "0000000000000000000000000000000000000000000000000000000000000000", -- 02
   "0000000000000000000000000000000000000000000000000000000000000000", -- 03
   "0000000000000000000000000000000000000000000000000000000000000000", -- 04
   "0000000000000000000000000000000000000000000000000000000000000000", -- 05
   "0000000000000000000000000000000000000000000000000000000000000000", -- 06
   "0000000000000000000000000000000000000000000000000000000000000000", -- 07
   "0000000000000000000000000000000000000000000000000000000000000000", -- 08
   "0000000000000000000000000000000000000000000000000000000000000000", -- 09
   "0000000000000000100000000000000000000000000000001000000000000000", -- 0a
   "0000000000000000100000000000000000000000000000001000000000000000", -- 0b
   "0000000000000111111000000000000000000000000001111110000000000000", -- 0c
   "0000000000001111111100000000000000000000000011111111000000000000", -- 0d
   "0000000000000111111000000000000000000000000001111110000000000000", -- 0e
   "0000000000000000100000000000000000000000000000001000000000000000", -- 0f
   "0000000000000000100000000000000000000000000000001000000000000000", -- 10
   "0000000000000000000000000000000000000000000000000000000000000000", -- 11
   "0000000000000000000000000000000000000000000000000000000000000000", -- 12
   "0000000000000000000000000000000000000000000000000000000000000000", -- 13
   "0000000000000000000000000000000000000000000000000000000000000000", -- 14
   "0000000000000000000000000000000000000000000000000000000000000000", -- 15
   "0000000000000000000000000000000000000000000000000000000000000000", -- 16
   "0000000000000000000000000000000000000000000000000000000000000000", -- 17
   "0000000000000000000000000000000000000000000000000000000000000000", -- 18
   "0000000000000000000000000000000000000000000000000000000000000000", -- 19
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1a
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1b
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1c
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1d
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1e
   "0000000000000000000000000000000000000000000000000000000000000000", -- 1f
   "0000000000000000000000000000000000000000000000000000000000000000", -- 20
   "0000000000000000000000000000000000000000000000000000000000000000", -- 21
   "0000000000000000000000000000000000000000000000000000000000000000", -- 22
   "0000000000000000000000000000000000000000000000000000000000000000", -- 23
   "0000000000000000000000000000000000000000000000000000000000000000", -- 24
   "0000000000000000000000000000000000000000000000000000000000000000", -- 25
   "0000000000000000000000000000000000000000000000000000000000000000", -- 26
   "0000000000000000000000000000000000000000000000000000000000000000", -- 27
   "0000000000000000000000000000000000000000000000000000000000000000", -- 28
   "0000000000000000000000000000000000000000000000000000000000000000", -- 29
   "0000000000000000100000000000000000000000000000001000000000000000", -- 2a
   "0000000000000000100000000000000000000000000000001000000000000000", -- 2b
   "0000000000000111111000000000000000000000000001111110000000000000", -- 2c
   "0000000000001111111100000000000000000000000011111111000000000000", -- 2d
   "0000000000000111111000000000000000000000000001111110000000000000", -- 2e
   "0000000000000000100000000000000000000000000000001000000000000000", -- 2f
   "0000000000000000100000000000000000000000000000001000000000000000", -- 30
   "0000000000000000000000000000000000000000000000000000000000000000", -- 31
   "0000000000000000000000000000000000000000000000000000000000000000", -- 32
   "0000000000000000000000000000000000000000000000000000000000000000", -- 33
   "0000000000000000000000000000000000000000000000000000000000000000", -- 34
   "0000000000000000000000000000000000000000000000000000000000000000", -- 35
   "0000000000000000000000000000000000000000000000000000000000000000", -- 36
   "0000000000000000000000000000000000000000000000000000000000000000", -- 37
   "0000000000000000000000000000000000000000000000000000000000000000", -- 38
   "0000000000000000000000000000000000000000000000000000000000000000", -- 39
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3a
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3b
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3c
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3d
   "0000000000000000000000000000000000000000000000000000000000000000", -- 3e
   "0000000000000000000000000000000000000000000000000000000000000000"  -- 3f
   );                            
      
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= ROM(to_integer(unsigned(addr_reg)));
end arch;
